-------------------------------------------------------------------------
-- Henry Duwe
-- Department of Electrical and Computer Engineering
-- Iowa State University
-------------------------------------------------------------------------


-- mux2t1_N.vhd
-------------------------------------------------------------------------
-- DESCRIPTION: This file contains an implementation of an N-bit wide 2:1
-- mux using structural VHDL, generics, and generate statements.
--
--
-- NOTES:
-- 1/6/20 by H3::Created.
-------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

entity addsub_n is
  generic(N : integer := 32); -- Generic of type integer for input/output data width. Default value is 32.
  port(nAdd_Sub    : in std_logic;
       i_A         : in std_logic_vector(N-1 downto 0);
       i_B         : in std_logic_vector(N-1 downto 0);
       o_S         : out std_logic_vector(N-1 downto 0);
       o_C         : out std_logic);

end addsub_n;

architecture structural of addsub_n is

  component adder_n is
	generic(N : integer := 32);
 	port(i_C          : in std_logic;
        i_X1         : in std_logic_vector(N-1 downto 0);
        i_X2         : in std_logic_vector(N-1 downto 0);
        o_S          : out std_logic_vector(N-1 downto 0);
        o_C          : out std_logic);
  end component;

  component mux2t1_n is
	generic(N : integer := 32);
  	port(i_S          : in std_logic;
        i_D0         : in std_logic_vector(N-1 downto 0);
        i_D1         : in std_logic_vector(N-1 downto 0);
        o_O          : out std_logic_vector(N-1 downto 0));
  end component;

  component onescomp_n is
	generic(N : integer := 32);
  	port(i_N         : in std_logic_vector(N-1 downto 0);
        o_O         : out std_logic_vector(N-1 downto 0));
  end component;
  signal start : std_logic_vector(N-1 downto 0);
  signal inverted : std_logic_vector(N-1 downto 0);

  signal temp : std_logic_vector(N-1 downto 0);
  signal muxOut : std_logic_vector(N-1 downto 0);
  signal final : std_logic_vector(N-1 downto 0);
  signal s_outC: std_logic;
begin

negation: process(s_outC, nAdd_Sub) is begin
  if nAdd_Sub = '1' then
	o_C <= not(s_outC);
  else
	o_C <= s_outC;
  end if;
end process negation;
  -- Instantiate N mux instances.
  G_NBit_ADDER: adder_n
  generic map(N => 32)
  port map(
              i_C      => nAdd_Sub,      -- All instances share the same select input.
              i_X1     => i_A,  -- ith instance's data 0 input hooked up to ith data 0 input.
              i_X2     => muxOut,  -- ith instance's data 1 input hooked up to ith data 1 input.
              o_S      => o_S,  -- ith instance's data output hooked up to ith data output.
	      o_C      => s_outC);

  G_NBit_MUX: mux2t1_n
  generic map(N => 32)
  port map(
              i_S      => nAdd_Sub,      -- All instances share the same select input.
              i_D0     => i_B,  -- ith instance's data 0 input hooked up to ith data 0 input.
              i_D1     => inverted,  -- ith instance's data 1 input hooked up to ith data 1 input.
              o_O      => muxOut);  -- ith instance's data output hooked up to ith data output.
 

  G_NBit_OCN: onescomp_n
  generic map(N => 32)
  port map(
              i_N     => i_B,  -- ith instance's data 0 input hooked up to ith data 0 input.
              o_O      => inverted);  -- ith instance's data output hooked up to ith data output.
  	  
end structural;
